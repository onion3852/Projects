module sram_controller (
    
);
    
endmodule