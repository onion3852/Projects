module tb_sram_controller();

endmodule